module motionestimator(
	input clk,
	input reset_n,
	output reg rdy,
	input en,
	// Inputs
	input  [9:0] ix,
	input  [9:0] iy,
	input  intra,    // Intra-coded macroblock, assume prediction = 128
	// Avalon Master
	output read,
	output write,
	output [31:0] addr,
	output [7:0]  writedata,
	input  [7:0]  readdata,
	input  waitrequest,
	input  readdatavalid,
	// Camera Interface
	output [9:0] x,
	output [9:0] y,
	output reg [1:0] cc,
	input  [7:0] px,
	// Output Interface
	input [7:0] raddr,
	output [15:0] q,
	input [7:0]  dctaddr,
	input [15:0] dctdata,
	output [9:0] xmin, // Motion vectors
	output [9:0] ymin);

	// Offsets generated by the block comparator
	wire [3:0] mx, my;
	// Address buses: waddr for writing the current macroblock to the MBRAM,
	// baddr for indexing into the camera's data
	wire [7:0] waddr, baddr;
	wire [15:0] wdata;
	// Current and old accumulator values
	wire [17:0] accum, oldaccum;
	reg  [17:0] next_accum;
	wire wren, mreq;
	reg cmp_en;

	// Current state
	wire [3:0] state;
	reg  [3:0] next_state;

	// Origin X, Y, and Offset DX, DY
	wire [9:0] ox, oy, dx, dy;
	reg [9:0] next_ox, next_oy, next_dx, next_dy;
	// Current search radius S
	wire [3:0] s;
	reg [3:0] next_s;
	// DX and DY values which produce the minimum value of accum
	wire [9:0] min_dx, min_dy;
	reg  [9:0] next_min_dx, next_min_dy;

	register #(18) ACCUM(.clk(clk), .in(reset_n  ? next_accum : 18'b0), .out(oldaccum), .en(1'b1));
	register #(10) OX(.clk(clk), .in(reset_n ? next_ox : 10'b0), .out(ox), .en(1'b1));
	register #(10) OY(.clk(clk), .in(reset_n ? next_oy : 10'b0), .out(oy), .en(1'b1));
	register #(10) DX(.clk(clk), .in(reset_n ? next_dx : 10'b0), .out(dx), .en(1'b1));
	register #(10) DY(.clk(clk), .in(reset_n ? next_dy : 10'b0), .out(dy), .en(1'b1));
	register #(10) MIN_DX(.clk(clk), .in(reset_n ? next_min_dx : 10'b0), .out(min_dx), .en(1'b1));
	register #(10) MIN_DY(.clk(clk), .in(reset_n ? next_min_dy : 10'b0), .out(min_dy), .en(1'b1));
	register #(4)  S(.clk(clk), .in(reset_n ? next_s : 4'b0), .out(s), .en(1'b1));
	register #(4)  STATE(.clk(clk), .in(reset_n ? next_state : 4'b0), .out(state), .en(1'b1));

	mbram external(.clock(clk), .data(wdata), .rdaddress(raddr),
		.wraddress(waddr), .wren(wren), .q(q));

	blkcompare comparator(.clk(clk), .reset_n(reset_n), .rdy(cmp_rdy), .en(cmp_en), .baddr(baddr),
		.bq(bq), .mx(mx), .my(my), .mq(intra ? 8'd128 : readdata), .mreq(mreq), .m_wait(intra ? 1'b0 : waitrequest), .m_valid(intra ? 1'b1 : readdatavalid),
		.waddr(waddr), .wdata(wdata), .wren(wren), .oldaccum(oldaccum), .accum(accum), .valid(valid));

	assign read = intra ? 1'b0 : mreq;

	assign x = ox + dx + baddr[3:0];
	assign y = oy + dy + baddr[7:4];
	
	always @(*) begin
		rdy = 1'b0;
		cc  = 2'b0;
		next_accum = oldaccum;
		next_ox = ox;
		next_oy = oy;
		next_dx = dx;
		next_dy = dy;
		next_min_dx = dx;
		next_min_dy = dy;
		next_s = s;
		next_state = state;
		case (state)
			4'h0: begin // Reset state
				rdy = 1'b1;
				if (en) begin
					next_ox = ix;
					next_oy = iy;
					next_dx = 10'b0;
					next_dy = 10'b0;
					next_min_dx = 10'b0;
					next_min_dy = 10'b0;
					next_s = 4'h4;
					next_accum = 18'h1FFFF;
					if (intra) begin
						next_state = 4'h1;
					end else begin
						next_state = 4'hF;
					end
				end
			end
			4'h1: begin // Intra compression start state
				if (cmp_rdy) begin
					next_state = 4'h2;
					cmp_en = 1'b1;
				end
			end
			4'h2: begin // Wait for the comparator to complete
				cc = 2'b00; // Select Y
				if (cmp_rdy) begin
					next_state = 4'h0;
				end
			end
			default: begin
				next_state = 4'h0;
			end
		endcase
	end
endmodule
