module motionestimator(
	input clk,
	input reset_n,
	output reg rdy,
	input en,
	input writeback, // If true, en signals writing back to Avalon
	// Inputs
	input  [9:0] ix,
	input  [9:0] iy,
	input  [31:0] base, // Avalon base address, for reading and writing
	input  intra,    // Intra-coded macroblock, assume prediction = 128
	// Avalon Master
	output read,
	output reg write,
	output [31:0] addr,
	output reg [7:0] writedata,
	input  [7:0]  readdata,
	input  waitrequest,
	input  readdatavalid,
	// Camera Interface
	output [9:0] x,
	output [9:0] y,
	output reg [1:0] cc,
	input  [7:0] px,
	// Motion vectors
	output [9:0] xmin,
	output [9:0] ymin,
	// Output Interface
	input [7:0] raddr,
	output [15:0] q,
	input [7:0]  dctaddr,
	input [15:0] dctdata,
	input dctwren
	);

	parameter WIDTH  = 10'd640;
	parameter HEIGHT = 10'd480;
	parameter YSIZE  = 32'd307200; // WIDTH * HEIGHT
	parameter UVSIZE = 32'd76800;  // WIDTH * HEIGHT / 4, for downsampling

	reg  [31:0] base_addr; // Base of current component
	// Offsets generated by the block comparator
	wire [3:0] mx, my, bx, by, wx, wy;
	// Address buses: waddr for writing the current macroblock to the MBRAM,
	// baddr for indexing into the camera's data
	wire [8:0]  waddr, baddr, dwaddr, draddr, paddr;
	wire [15:0] wdata, pq, bq, data;
	// Current and old accumulator values
	wire [17:0] accum, oldaccum;
	reg  [17:0] next_accum;
	wire wren, mreq, cmp_rdy, valid;
	reg cmp_en, wsel, dsel;

	// Current state
	wire [3:0] state;
	reg  [3:0] next_state;
	
	wire [1:0] bcc, wcc;
	reg  [1:0] next_cc;

	// Origin X, Y, and Offset DX, DY
	wire [9:0] ox, oy, dx, dy;
	reg [9:0] next_ox, next_oy, next_dx, next_dy;
	// Current search radius S
	wire [3:0] s, min_s;
	reg [3:0] next_s, next_min_s;
	// Next values for the motion vectors
	wire [9:0] min_dx, min_dy;
	reg  [9:0] next_min_dx, next_min_dy;
	
	wire [3:0] max;
	reg  [3:0] next_max;

	register #(18) ACCUM(.clk(clk), .in(reset_n  ? next_accum : 18'b0), .out(oldaccum), .en(1'b1));
	register #(10) OX(.clk(clk), .in(reset_n ? next_ox : 10'b0), .out(ox), .en(1'b1));
	register #(10) OY(.clk(clk), .in(reset_n ? next_oy : 10'b0), .out(oy), .en(1'b1));
	register #(10) DX(.clk(clk), .in(reset_n ? next_dx : 10'b0), .out(dx), .en(1'b1));
	register #(10) DY(.clk(clk), .in(reset_n ? next_dy : 10'b0), .out(dy), .en(1'b1));
	register #(10) MIN_DX(.clk(clk), .in(reset_n ? next_min_dx : 10'b0), .out(min_dx), .en(1'b1));
	register #(10) MIN_DY(.clk(clk), .in(reset_n ? next_min_dy : 10'b0), .out(min_dy), .en(1'b1));
	register #(4)  S(.clk(clk), .in(reset_n ? next_s : 4'b0), .out(s), .en(1'b1));
	register #(4)  MIN_S(.clk(clk), .in(reset_n ? next_min_s : 4'b0), .out(min_s), .en(1'b1));
	register #(4)  STATE(.clk(clk), .in(reset_n ? next_state : 4'b0), .out(state), .en(1'b1));
	register #(2)  CC(.clk(clk), .in(reset_n ? next_cc : 2'b0), .out(wcc), .en(1'b1));
	register #(4)  MAX(.clk(clk), .in(reset_n ? next_max : 4'b0), .out(max), .en(1'b1));

	mbram predicted(.clock(clk), .data(intra ? 16'd128 : {8'b0, readdata}), .rdaddress(paddr),
		.wraddress(waddr), .wren(wren), .q(pq));

	mbram external(.clock(clk), .data(wdata), .rdaddress(wsel ? paddr : (dsel ? draddr : baddr)),
		.wraddress(dwaddr), .wren(wren), .q(q));

	blkcompare comparator(.clk(clk), .reset_n(reset_n), .rdy(cmp_rdy), .en(cmp_en), .cc(bcc), .bx(bx), .by(by),
		.bq(bq), .mx(mx), .my(my), .mq(intra ? 8'd128 : readdata), .mreq(mreq), .m_wait(intra ? 1'b0 : waitrequest), .m_valid(intra ? 1'b1 : readdatavalid),
		.wx(wx), .wy(wy), .wdata(wdata), .wren(wren), .oldaccum(oldaccum), .accum(accum), .valid(valid));

	XYCCtoAddr BADDR(.x(bx), .y(by), .cc(cc), .addr(baddr));
	XYCCtoAddr WADDR(.x(wx), .y(wy), .cc(cc), .addr(waddr));
	XYCCtoAddr DCTWADDR(.x(dctaddr[3:0]), .y(dctaddr[7:4]), .cc(cc), .addr(dwaddr));
	XYCCtoAddr DCTRADDR(.x(raddr[3:0]), .y(raddr[7:4]), .cc(cc), .addr(draddr));
	XYCCtoAddr PADDR(.x(dx[3:0]), .y(dy[3:0]), .cc(cc), .addr(paddr));

	assign read = intra ? 1'b0 : mreq;
	assign x = ox + dx + bx;
	assign y = oy + dy + by;
	assign xmin = (ox - ix) + min_dx;
	assign ymin = (oy - iy) + min_dy;
	assign data = pq + q;
	assign addr = base_addr + (wsel ? iy + dy : y) * WIDTH + (wsel ? ix + dx : x);
	
	always @(*) begin
		case (cc)
			2'b00: begin
				base_addr = base;
			end
			2'b01: begin
				base_addr = base + YSIZE;
			end
			2'b10: begin
				base_addr = base + YSIZE + UVSIZE;
			end
			default: begin
				base_addr = 32'b0;
			end
		endcase
	end

	always @(*) begin
		rdy = 1'b0;
		write = 1'b0;
		wsel = 1'b0;
		dsel = 1'b0;
		next_accum = oldaccum;
		next_ox = ox;
		next_oy = oy;
		next_dx = dx;
		next_dy = dy;
		next_min_dx = dx;
		next_min_dy = dy;
		next_max = max;
		next_s = s;
		next_min_s = min_s;
		next_state = state;
		next_cc = wcc;
		cc = bcc;
		case (state)
			4'h0: begin // Reset state
				rdy = 1'b1;
				dsel = 1'b1;
				if (en) begin
					next_ox = ix;
					next_oy = iy;
					next_dx = 10'b0;
					next_dy = 10'b0;
					next_min_dx = 10'b0;
					next_min_dy = 10'b0;
					next_s = 4'h4;
					next_accum = 18'h1FFFF;
					next_cc = 2'b0;
					if (writeback) begin
						next_state = 4'h5;
					end else begin
						if (intra) begin
							next_state = 4'h1;
						end else begin
							next_state = 4'h3;
						end
					end
				end
			end
			4'h1: begin // Intra compression start state
				if (cmp_rdy) begin
					next_state = 4'h2;
					cmp_en = 1'b1;
				end
			end
			4'h2: begin // Wait for the comparator to complete
				if (cmp_rdy) begin
					next_state = 4'h0;
				end
			end
			4'h3: begin // Inter compression start state
				if (cmp_rdy) begin
					cmp_en = 1'b1;
					if (($signed(ox - dx) < $signed(10'd0))
					|| (ox > (WIDTH - 10'd16))
					|| (oy > (HEIGHT - 10'd16))
					|| ($signed(oy - dy) < $signed(10'd0)))
					 begin
						// Clipping: Entire macroblock must be within image
						cmp_en = 1'b0;
					end
					next_state = 4'h4;
				end
			end
			4'h4: begin // Inter compression wait state
				if (cmp_rdy) begin
					if (valid) begin
						next_accum = accum;
						next_min_dx = dx;
						next_min_dy = dy;
						next_min_s = s;
					end
					if ((dx == 10'd0) && (dy == 10'd0)) begin
						next_dy = 10'd0 - {6'd0,s};
					end else if ((dx == 10'd0) && (dy == (10'd0 - {6'd0,s}))) begin
						next_dx = {6'd0,s};
					end else if ((dx == {6'd0,s}) && (dy == (10'd0 - {6'd0,s}))) begin
						next_dy = 10'd0;
					end else if ((dx == {6'd0,s}) && (dy == 10'd0)) begin
						next_dy = {6'd0,s};
					end else if ((dx == {6'd0,s}) && (dy == {6'd0,s})) begin
						next_dx = 10'd0;
					end else if ((dx == 10'd0) && (dy == {6'd0, s})) begin
						next_dx = 10'd0 - {6'd0,s};
					end else if ((dx == 10'd0 - {6'd0,s}) && (dy == {6'd0,s})) begin
						next_dy = 10'd0;
					end else if ((dx == 10'd0 - {6'd0,s}) && (dy == 10'd0)) begin
						next_dy = 10'd0 - {6'd0,s};
					end else begin
						// After checking S = 0 and S = 4, continue to S = 1
						if (s == 4'd4) begin
							next_s = 4'd1;
						// Then, if the minimum occurs at S = 0, exit
						end else if (min_s == 4'd0) begin
							next_state = 4'h0;
						// Else if S = 1, restart from S = 1 and then exit
						end else if (s == 4'd1) begin
							if ((ox == ix) && (oy == iy)) begin
								next_ox = ox + min_dx;
								next_oy = oy + min_dy;
								next_dx = 10'd0;
								next_dy = -10'd1;
							end else begin
								next_state = 4'h0;
							end
						end else begin // min_s == 4 or 2
							next_ox = ox + min_dx;
							next_oy = oy + min_dy;
							next_dx = 10'd0;
							next_dy = 10'd0 - {7'd0,s[3:1]};
							next_s  = {1'd0, s[3:1]};
						end
					end
				end
			end
			4'h5: begin // Write YUV back to Avalon
				cc = wcc;
				wsel = 1'b1;
				if ($signed(data) < 16'd0) begin
					writedata = 8'd0;
				end else if ($signed(data) > 16'd255) begin
					writedata = 8'd255;
				end else begin
					writedata = data[7:0];
				end
				if (!waitrequest) begin
					write = 1'b1;
					next_dx = dx + 4'h1;
					if (dx == max) begin
						if (dy == max) begin
							next_cc = wcc + 2'b01;
							next_max = 4'd7;
							if (cc == 2'b10) begin
								next_state = 4'h0;
							end
							next_dx = max;
						end else begin
							next_dx = 4'd0;
							next_dy = dy + 4'd1;
						end
					end

				end
			end
			default: begin
				next_state = 4'h0;
			end
		endcase
	end
endmodule
